file1 add klajsdlakdj

